`define NOP   4'b0000
`define STORE 4'b0001
`define LOAD  4'b0010
`define ADDC  4'b0011
`define SUBC  4'b0100
`define AND   4'b0101
`define OR    4'b0110
`define XOR   4'b0111
`define SHL   4'b1000
`define SHR   4'b1001
`define SHRA  4'b1010
`define ADDI  4'b1011
`define SUBI  4'b1100
`define ANDI  4'b1101
`define ORI   4'b1110
`define XORI  4'b1111